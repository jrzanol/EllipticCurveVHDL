LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

PACKAGE MYWORK IS

-- Definições da Curva Elíptica: https://github.com/vjudeu/curves1000/blob/master/bits/bits64.txt
CONSTANT P : STD_LOGIC_VECTOR (63 DOWNTO 0) := X"fffffffefffff833"; -- Primo
CONSTANT Gx : STD_LOGIC_VECTOR (63 DOWNTO 0) := X"90fab331bd548cce"; -- Pk=1
CONSTANT Gy : STD_LOGIC_VECTOR (63 DOWNTO 0) := X"1d8f41753fd04b4a";
CONSTANT Gx2 : STD_LOGIC_VECTOR (63 DOWNTO 0) := X"f7e97ff3a83de0e3"; -- Pk=2
CONSTANT Gy2 : STD_LOGIC_VECTOR (63 DOWNTO 0) := X"9023999ee95d53d3";

COMPONENT AddOnePoint IS
PORT(CLK, RST, START: IN STD_LOGIC;
		X1, Y1: IN SIGNED (63 DOWNTO 0);
		XOUT, YOUT: OUT SIGNED (63 DOWNTO 0);
		DONE: OUT STD_LOGIC);
END COMPONENT;

COMPONENT ModAdd IS
PORT(X1, X2: IN SIGNED (63 DOWNTO 0);
		XOUT: OUT SIGNED (63 DOWNTO 0));
END COMPONENT;

COMPONENT ModSub IS
PORT(X1, X2: IN SIGNED (63 DOWNTO 0);
		XOUT: OUT SIGNED (63 DOWNTO 0));
END COMPONENT;

COMPONENT ModMult IS
PORT(A, B: IN SIGNED(63 DOWNTO 0);
		XOUT: OUT SIGNED(63 DOWNTO 0));
END COMPONENT;

COMPONENT ModNeg IS
PORT(X1: IN SIGNED (63 DOWNTO 0);
		XOUT: OUT SIGNED (63 DOWNTO 0));
END COMPONENT;

COMPONENT ModInv IS
PORT(CLK, RESET, START: IN STD_LOGIC;
		A, B: IN UNSIGNED(63 downto 0);
		DONE: OUT STD_LOGIC;
		INVERSE: OUT UNSIGNED(63 downto 0));
END COMPONENT;

END PACKAGE;

